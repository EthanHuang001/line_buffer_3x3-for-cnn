module window_3x3 #(
    parameter DATA_WIDTH = 8,
    parameter WIDTH      = 640,
    parameter HEIGHT     = 480
)(
    input  wire                   clk,
    input  wire                   rst_n,
    
    input  wire                   in_valid,     // ������"����"��Ч
    input  wire [DATA_WIDTH-1:0]  pix_curr,     // ��ǰ�� y
    input  wire [DATA_WIDTH-1:0]  pix_m1,       // y-1 ��
    input  wire [DATA_WIDTH-1:0]  pix_m2,       // y-2 ��
    
    output reg                   win_valid,    // 3x3 ������Ч
    output wire [DATA_WIDTH-1:0]  p00, p01, p02,
    output wire [DATA_WIDTH-1:0]  p10, p11, p12,
    output wire [DATA_WIDTH-1:0]  p20, p21, p22
);

// �ڲ��Ĵ�������
reg [DATA_WIDTH-1:0] p00_reg, p01_reg, p02_reg;
reg [DATA_WIDTH-1:0] p10_reg, p11_reg, p12_reg;
reg [DATA_WIDTH-1:0] p20_reg, p21_reg, p22_reg;

// ������Ч��־�Ĵ���
reg win_valid_reg;
// ��������ѡ����
wire [DATA_WIDTH-1:0] pix_m2_in = in_valid ? pix_m2 : {DATA_WIDTH{1'b0}};
wire [DATA_WIDTH-1:0] pix_m1_in = in_valid ? pix_m1 : {DATA_WIDTH{1'b0}};
wire [DATA_WIDTH-1:0] pix_curr_in = in_valid ? pix_curr : {DATA_WIDTH{1'b0}};

// ����λ�߼�
always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        // ��λ���мĴ���
        p00_reg <= {DATA_WIDTH{1'b0}};
        p01_reg <= {DATA_WIDTH{1'b0}};
        p02_reg <= {DATA_WIDTH{1'b0}};
        
        p10_reg <= {DATA_WIDTH{1'b0}};
        p11_reg <= {DATA_WIDTH{1'b0}};
        p12_reg <= {DATA_WIDTH{1'b0}};
        
        p20_reg <= {DATA_WIDTH{1'b0}};
        p21_reg <= {DATA_WIDTH{1'b0}};
        p22_reg <= {DATA_WIDTH{1'b0}};
        
        win_valid_reg <= 1'b0;
    end
    else begin
        // ��һ����λ: pix_m2
        p02_reg <= p01_reg;  // p01 -> p02
        p01_reg <= p00_reg;  // p00 -> p01
        p00_reg <= pix_m2_in; // ������ -> p00
        
        // �ڶ�����λ: pix_m1
        p12_reg <= p11_reg;  // p11 -> p12
        p11_reg <= p10_reg;  // p10 -> p11
        p10_reg <= pix_m1_in; // ������ -> p10
        
        // ��������λ: pix_curr
        p22_reg <= p21_reg;  // p21 -> p22
        p21_reg <= p20_reg;  // p20 -> p21
        p20_reg <= pix_curr_in; // ������ -> p20
        
        // ������Ч�ź�����
        // �����������2����Ч��ʱ�����ڿ�ʼ��Ч
        win_valid_reg <= in_valid;
		win_valid <= win_valid_reg;
    end
end

// �������
assign p02 = p00_reg;
assign p01 = p01_reg;
assign p00 = p02_reg;
assign p12 = p10_reg;
assign p11 = p11_reg;
assign p10 = p12_reg;
assign p22 = p20_reg;
assign p21 = p21_reg;
assign p20 = p22_reg;

endmodule