`timescale 1ns / 1ps

module line_buffer_3x3 #(
    parameter DATA_WIDTH = 8,
    parameter WIDTH      = 640,   // һ�������� (<=1024)
    parameter HEIGHT     = 480    // ͼ��߶ȣ���ʵ������
)(
    input  wire                   clk,
    input  wire                   rst_n,

    input  wire                   in_valid,     // ����������Ч
    input  wire [DATA_WIDTH-1:0]  pix_in,       // ��ͨ����������

    // ����� window_3x3 �� 3x3 ����
    output wire                   win_valid,
    output wire [DATA_WIDTH-1:0]  p00, p01, p02,
    output wire [DATA_WIDTH-1:0]  p10, p11, p12,
    output wire [DATA_WIDTH-1:0]  p20, p21, p22
);

    // ======================================================
    // 1) ��/�м��������� in_valid ��������ʵ��������У�
    // ======================================================
    reg [9:0]   x_cnt;   // �м���
    reg [15:0]  y_cnt;   // �м��� (0..HEIGHT-1)

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            x_cnt <= 10'd0;
            y_cnt <= 16'd0;
        end else if (in_valid) begin
            if (x_cnt == WIDTH-1) begin
                x_cnt <= 10'd0;
                if (y_cnt < HEIGHT-1)
                    y_cnt <= y_cnt + 1'b1;
            end else begin
                x_cnt <= x_cnt + 1'b1;
            end
        end
    end

    // ======================================================
    // 2) ������ˮ�������ĸ� window
    //    ����pix_curr_s1_stream / y_cnt_d2 / x_cnt_d2 / in_v_d2
    // ======================================================
    reg                  in_v_d1, in_v_d2;
    reg [9:0]            x_cnt_d1, x_cnt_d2;
    reg [15:0]           y_cnt_d1, y_cnt_d2;
    reg [DATA_WIDTH-1:0] pix_d1;
    reg [DATA_WIDTH-1:0] pix_curr_s1_stream;   // ������ģʽ���¸� window �ĵ�ǰ������

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            in_v_d1            <= 1'b0;
            in_v_d2            <= 1'b0;
            x_cnt_d1           <= 10'd0;
            x_cnt_d2           <= 10'd0;
            y_cnt_d1           <= 16'd0;
            y_cnt_d2           <= 16'd0;
            pix_d1             <= {DATA_WIDTH{1'b0}};
            pix_curr_s1_stream <= {DATA_WIDTH{1'b0}};
        end else begin
            // ��һ��
            in_v_d1 <= in_valid;
            if (in_valid) begin
                x_cnt_d1 <= x_cnt;
                y_cnt_d1 <= y_cnt;
                pix_d1   <= pix_in;
            end

            // �ڶ���
            in_v_d2 <= in_v_d1;
            if (in_v_d1) begin
                x_cnt_d2           <= x_cnt_d1;
                y_cnt_d2           <= y_cnt_d1;
                pix_curr_s1_stream <= pix_d1;
            end
        end
    end

    // ======================================================
    // 3) �ײ� padding ���ƣ������һ����Ч���ݽ������ BOTTOM_GAP �ģ������һ��
    // ======================================================
    localparam BOTTOM_GAP = 5;

    reg        padding_mode;      // 1����������� padding ��
    reg [2:0]  gap_cnt;           // �հ׼���
    reg [9:0]  bottom_x_cnt;      // ����ɨ���� (0..WIDTH)
    reg        frame_done_pulse;  // һ֡�������壨������� RAM��

    wire last_pixel_2nd_stage;
    assign last_pixel_2nd_stage =
        in_v_d2 &&
        (y_cnt_d2 == (HEIGHT-1)) &&
        (x_cnt_d2 == (WIDTH-1));

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            padding_mode     <= 1'b0;
            gap_cnt          <= 3'd0;
            bottom_x_cnt     <= 10'd0;
            frame_done_pulse <= 1'b0;
        end else begin
            frame_done_pulse <= 1'b0;   // Ĭ������

            if (!padding_mode) begin
                // ����ģʽ���ȴ����һ�����ؽ���ڶ���
                if (last_pixel_2nd_stage) begin
                    gap_cnt <= 3'd1;
                end else if (gap_cnt != 3'd0 && gap_cnt < BOTTOM_GAP) begin
                    gap_cnt <= gap_cnt + 1'b1;
                end else if (gap_cnt == BOTTOM_GAP) begin
                    // GAP ���������� padding ��
                    padding_mode <= 1'b1;
                    bottom_x_cnt <= 10'd0;
                    gap_cnt      <= 3'd0;
                end
            end else begin
                // padding_mode: bottom_x_cnt �� 0 ���� WIDTH
                if (bottom_x_cnt == WIDTH) begin
                    // ��һ�ģ������һ�����ص� q ����ˮ�������ʱ��
                    padding_mode     <= 1'b0;
                    bottom_x_cnt     <= 10'd0;
                    frame_done_pulse <= 1'b1;   // �� һ֡�������� RAM
                end else begin
                    bottom_x_cnt <= bottom_x_cnt + 1'b1;
                end
            end
        end
    end

    // �� RAM �Ķ���ַ & ��ʹ��
    wire [9:0] addr_x_for_ram = padding_mode ? bottom_x_cnt : x_cnt;
    wire       rden_for_ram   = padding_mode ? (bottom_x_cnt < WIDTH) : in_valid;

    // ======================================================
    // 4) ������ RAM���� aclr �� register IP
    // ======================================================
    wire [9:0] ram0_rdaddr = addr_x_for_ram;
    wire [9:0] ram1_rdaddr = addr_x_for_ram;
    wire       ram0_rden   = rden_for_ram;
    wire       ram1_rden   = rden_for_ram;

    reg  [DATA_WIDTH-1:0] ram0_data;
    reg  [9:0]            ram0_wraddr;
    reg                   ram0_wren;
    wire [DATA_WIDTH-1:0] ram0_q;

    reg  [DATA_WIDTH-1:0] ram1_data;
    reg  [9:0]            ram1_wraddr;
    reg                   ram1_wren;
    wire [DATA_WIDTH-1:0] ram1_q;

    // ��� IP��
    // register(aclr, clock, data, rdaddress, wraddress, wren, rden, q);
    register u_ram0 (
        .aclr     (frame_done_pulse),  // �� һ֡����ʱ�첽����
        .clock    (clk),
        .data     (ram0_data),
        .rdaddress(ram0_rdaddr),
        .wraddress(ram0_wraddr),
        .wren     (ram0_wren),
        .rden     (ram0_rden),
        .q        (ram0_q)
    );

    register u_ram1 (
        .aclr     (frame_done_pulse),  // �� һ֡����ʱ�첽����
        .clock    (clk),
        .data     (ram1_data),
        .rdaddress(ram1_rdaddr),
        .wraddress(ram1_wraddr),
        .wren     (ram1_wren),
        .rden     (ram1_rden),
        .q        (ram1_q)
    );

    // ======================================================
    // 5) ��ֱ 3 ���� & д��ƹ��
    // ======================================================
    // padding ��ʹ�������к� HEIGHT����ʵֻӰ�� m1/m2 ��ѡ��
    wire [15:0] y_for_window = padding_mode ? HEIGHT[15:0] : y_cnt_d2;

    // �����͸� window �� curr
    wire [DATA_WIDTH-1:0] pix_curr_s1 =
        padding_mode           ? {DATA_WIDTH{1'b0}} :   // ���� curr = 0
        (in_v_d2              ) ? pix_curr_s1_stream :
                                  {DATA_WIDTH{1'b0}};

    // m1/m2 �������
    wire [DATA_WIDTH-1:0] pix_m1_normal;
    wire [DATA_WIDTH-1:0] pix_m2_normal;

    assign pix_m1_normal =
        (y_for_window == 16'd0) ? {DATA_WIDTH{1'b0}} :           // ��������һ��
        (y_for_window == 16'd1) ? ram0_q :                       // ��1�е���һ���� RAM0
        ( ((y_for_window - 1) & 16'h0001) ? ram1_q : ram0_q );   // y-1�� -> RAM1, ż -> RAM0

    assign pix_m2_normal =
        (y_for_window <= 16'd1) ? {DATA_WIDTH{1'b0}} :           // ǰ������ y-2
        ( ((y_for_window - 2) & 16'h0001) ? ram1_q : ram0_q );   // y-2 ��ż�ж�

    // m1/m2 padding �У�m1 �����һ�У�m2 �õ����ڶ��У����ߵ���
    localparam [15:0] LAST_ROW = HEIGHT-1;

    wire last_row_is_odd  = LAST_ROW[0];   // 1: ���һ���к�Ϊ����
    wire [DATA_WIDTH-1:0] pix_m1_bottom =
        last_row_is_odd ? ram1_q : ram0_q; // m1 = ���һ��
    wire [DATA_WIDTH-1:0] pix_m2_bottom =
        last_row_is_odd ? ram0_q : ram1_q; // m2 = �����ڶ��У�ȡ����

    wire [DATA_WIDTH-1:0] pix_m1_s1 = padding_mode ? pix_m1_bottom : pix_m1_normal;
    wire [DATA_WIDTH-1:0] pix_m2_s1 = padding_mode ? pix_m2_bottom : pix_m2_normal;

    // д��ǰ�н� RAM��ƹ�ң�����ֻ������ģʽ��padding ģʽ��д
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            ram0_wraddr <= 10'd0;
            ram1_wraddr <= 10'd0;
            ram0_wren   <= 1'b0;
            ram1_wren   <= 1'b0;
            ram0_data   <= {DATA_WIDTH{1'b0}};
            ram1_data   <= {DATA_WIDTH{1'b0}};
        end else begin
            ram0_wren <= 1'b0;
            ram1_wren <= 1'b0;

            if (!padding_mode && in_v_d2) begin
                if (y_cnt_d2[0] == 1'b0) begin
                    // ż����д RAM0
                    ram0_wraddr <= x_cnt_d2;
                    ram0_data   <= pix_curr_s1_stream;
                    ram0_wren   <= 1'b1;
                end else begin
                    // ������д RAM1
                    ram1_wraddr <= x_cnt_d2;
                    ram1_data   <= pix_curr_s1_stream;
                    ram1_wren   <= 1'b1;
                end
            end
        end
    end

    // ======================================================
    // 6) �� window �� in_valid��
    //    �����У��ӵڶ��п�ʼ���������ֻ�� padding �����У�
    //    padding �У�bottom_valid_raw���������ӳ�һ�Ķ��� ram_q
    // ======================================================
    wire win_in_valid_normal = in_v_d2 && (y_cnt_d2 >= 16'd1);

    // padding �У�bottom_x_cnt = 0..WIDTH
    wire bottom_valid_raw = padding_mode && (bottom_x_cnt > 0) && (bottom_x_cnt <= WIDTH);

    // Ϊ�˺� RAM �� q ���룬padding ��Ч�ٴ�һ��
    reg bottom_valid_d1;
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n)
            bottom_valid_d1 <= 1'b0;
        else
            bottom_valid_d1 <= bottom_valid_raw;
    end

    wire win_in_valid = padding_mode ? bottom_valid_d1
                                     : win_in_valid_normal;

    // ======================================================
    // 7) window_3x3��������� shift + ���� padding
    // ======================================================
    window_3x3 #(
        .DATA_WIDTH(DATA_WIDTH),
        .WIDTH     (WIDTH),
        .HEIGHT    (HEIGHT)
    ) u_window_3x3 (
        .clk      (clk),
        .rst_n    (rst_n),
        .in_valid (win_in_valid),
        .pix_curr (pix_curr_s1),
        .pix_m1   (pix_m1_s1),
        .pix_m2   (pix_m2_s1),
        .win_valid(win_valid),
        .p00      (p00),
        .p01      (p01),
        .p02      (p02),
        .p10      (p10),
        .p11      (p11),
        .p12      (p12),
        .p20      (p20),
        .p21      (p21),
        .p22      (p22)
    );

endmodule
