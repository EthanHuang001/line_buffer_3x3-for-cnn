`timescale 1ns/1ps

module tb_window_3x3();

// ��������
parameter DATA_WIDTH = 8;
parameter CLK_PERIOD = 40;  // 100MHz
parameter WIDTH = 10;       // �򻯲��ԣ�ʹ�ý�С���
parameter HEIGHT = 8;

// �ź�����
reg clk;
reg rst_n;
reg in_valid;
reg [DATA_WIDTH-1:0] pix_curr;
reg [DATA_WIDTH-1:0] pix_m1;
reg [DATA_WIDTH-1:0] pix_m2;

wire win_valid;
wire [DATA_WIDTH-1:0] p00, p01, p02;
wire [DATA_WIDTH-1:0] p10, p11, p12;
wire [DATA_WIDTH-1:0] p20, p21, p22;

// ʱ������
always #(CLK_PERIOD/2) clk = ~clk;

// ʵ��������ģ��
window_3x3 #(
    .DATA_WIDTH(DATA_WIDTH),
    .WIDTH(WIDTH),
    .HEIGHT(HEIGHT)
) u_window_3x3 (
    .clk(clk),
    .rst_n(rst_n),
    .in_valid(in_valid),
    .pix_curr(pix_curr),
    .pix_m1(pix_m1),
    .pix_m2(pix_m2),
    .win_valid(win_valid),
    .p00(p00),
    .p01(p01),
    .p02(p02),
    .p10(p10),
    .p11(p11),
    .p12(p12),
    .p20(p20),
    .p21(p21),
    .p22(p22)
);

// ���Լ���
integer i, j;
integer pixel_value = 1;
integer clock_count = 0;

initial begin
    // ��ʼ��
    clk = 0;
    rst_n = 0;
    in_valid = 0;
    pix_curr = 0;
    pix_m1 = 0;
    pix_m2 = 0;
    pixel_value = 1;
    clock_count = 0;
    
    // ��λ
    #(CLK_PERIOD*2);
    rst_n = 1;
    
    $display("=========================================");
    $display("��ʼ���� 3x3 ����ģ��");
    $display("=========================================\n");
    
    // ����1: ����������
    $display("����1: ��������������");
    $display("ʱ������  in_valid ����ֵ(m2,m1,curr) ������Ч ��������");
    $display("-----------------------------------------------------------------");
    #(CLK_PERIOD/2);
    in_valid = 1;
    for (i = 0; i < 12; i = i + 1) begin
        pix_m2 = pixel_value;      // ��y-2
        pix_m1 = pixel_value + 1;  // ��y-1
        pix_curr = pixel_value + 2; // ��y
        
        #CLK_PERIOD;
        clock_count = clock_count + 1;
        
        // ��ʾ����״̬
        if (win_valid) begin
            $display("����%2d:  %8b  (%3d,%3d,%3d)    %8b  (%3d,%3d,%3d)", 
                    clock_count, in_valid, pix_m2, pix_m1, pix_curr, win_valid,
                    p00, p01, p02);
            $display("                       p10,p11,p12: (%3d,%3d,%3d)", 
                    p10, p11, p12);
            $display("                       p20,p21,p22: (%3d,%3d,%3d)", 
                    p20, p21, p22);
        end
        else begin
            $display("����%2d:  %8b  (%3d,%3d,%3d)    %8b  (�ȴ��������...)", 
                    clock_count, in_valid, pix_m2, pix_m1, pix_curr, win_valid);
        end
        
        pixel_value = pixel_value + 3;
    end
    
    // ����2: ģ��padding��in_valid=0����������λ��
    $display("\n����2: ģ��padding��in_valid=0��");
    $display("ʱ������  in_valid ����ֵ(m2,m1,curr) ������Ч ��������");
    $display("-----------------------------------------------------------------");
    
    in_valid = 0;
    for (i = 0; i < 5; i = i + 1) begin
        #CLK_PERIOD;
        clock_count = clock_count + 1;
        
        if (win_valid) begin
            $display("����%2d:  %8b  (%3d,%3d,%3d)    %8b  (%3d,%3d,%3d)", 
                    clock_count, in_valid, 0, 0, 0, win_valid,
                    p00, p01, p02);
            $display("                       p10,p11,p12: (%3d,%3d,%3d)", 
                    p10, p11, p12);
            $display("                       p20,p21,p22: (%3d,%3d,%3d)", 
                    p20, p21, p22);
        end
    end
    
    // ����3: ���¿�ʼ������
    $display("\n����3: ���¿�ʼ������");
    $display("ʱ������  in_valid ����ֵ(m2,m1,curr) ������Ч ��������");
    $display("-----------------------------------------------------------------");
    
    in_valid = 1;
    for (i = 0; i < 8; i = i + 1) begin
        pix_m2 = 100 + i*3;        // ��y-2
        pix_m1 = 101 + i*3;        // ��y-1
        pix_curr = 102 + i*3;      // ��y
        
        #CLK_PERIOD;
        clock_count = clock_count + 1;
        
        if (win_valid) begin
            $display("����%2d:  %8b  (%3d,%3d,%3d)    %8b  (%3d,%3d,%3d)", 
                    clock_count, in_valid, pix_m2, pix_m1, pix_curr, win_valid,
                    p00, p01, p02);
            $display("                       p10,p11,p12: (%3d,%3d,%3d)", 
                    p10, p11, p12);
            $display("                       p20,p21,p22: (%3d,%3d,%3d)", 
                    p20, p21, p22);
        end
    end
    
    // ��������
    #(CLK_PERIOD*5);
    $display("\n=========================================");
    $display("�������");
    $display("=========================================");
    $finish;
end

// ��ش��ڱ仯
always @(posedge clk) begin
    if (rst_n) begin
        if (win_valid) begin
            // ��������Ҫʱ��Ӹ���ϸ�ļ��
        end
    end
end

// ���沨���ļ�
initial begin
    $dumpfile("window_3x3.vcd");
    $dumpvars(0, tb_window_3x3);
end

endmodule